library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use ieee.math_real.all;

-- Include the package where the matrix is defined
use work.MatrixPkg.ALL;         -- Include the package with the matrix definition

entity FPGA_Edge_Detection is
    port (
        clk : in STD_LOGIC;             -- Clock input
        reset : in STD_LOGIC;           -- Reset input
        input_signal : in STD_LOGIC_VECTOR(7 downto 0);  -- Input signal
        segmentsL_i0 : out STD_LOGIC_VECTOR(6 downto 0);  -- 7-segment for i0
        segmentsL_i1 : out STD_LOGIC_VECTOR(6 downto 0);  -- 7-segment for i1
        segmentsL_i2 : out STD_LOGIC_VECTOR(6 downto 0);  -- 7-segment for i2
        segmentsL_i3 : out STD_LOGIC_VECTOR(6 downto 0)   -- 7-segment for i3
    );
end FPGA_Edge_Detection;

architecture STRUCT of FPGA_Edge_Detection is

    -- Matrix and filter variables from MatrixPkg
    signal processed_signal : STD_LOGIC_VECTOR(7 downto 0);
    signal edge_matrix : ImageMatrix;
    
    -- BCD signals for the 7-segment display
    signal i0_signal, i1_signal, i2_signal, i3_signal : STD_LOGIC_VECTOR(3 downto 0); -- BCD signals

    -- Function to compute the threshold value (mean of the matrix)
    function compute_threshold(my_matrix: ImageMatrix) return integer is
        variable sum : integer := 0;
        variable mean : integer := 1;
    begin
        -- Sum all the values in the image matrix
        for i in 0 to 9 loop 
            for j in 0 to 9 loop
                sum := sum + my_matrix(i, j);  -- Assuming my_matrix contains the image data
            end loop;
        end loop;

        -- Compute the mean (threshold)
        mean := sum / 100;  -- Assuming a 10x10 matrix (100 elements in total)
        return mean;
    end function;

    -- Function to compute gradient magnitude
    function compute_edge(x: integer; y: integer; T: integer) return integer is
        variable gx_val : integer := 0;
        variable gy_val : integer := 0;
        variable edge_val : integer := 0;
    begin
        for i in 0 to 2 loop
            for j in 0 to 2 loop
                -- Apply the Prewitt Gx and Gy filters on the image matrix
                gx_val := gx_val + (my_matrix(x+i, y+j) * Gx(i, j));
                gy_val := gy_val + (my_matrix(x+i, y+j) * Gy(i, j));
            end loop;
        end loop;

        -- Compute the magnitude of the gradient
        edge_val := integer(sqrt(real(gx_val**2 + gy_val**2)));

        -- Return edge based on threshold
        if edge_val < T then 
            return 0;
        else 
            return 1;
        end if;
    end function;

    -- Convert integer to STD_LOGIC_VECTOR (4 bits for BCD representation)
    function int_to_bcd(val : integer) return STD_LOGIC_VECTOR is
    begin
        return STD_LOGIC_VECTOR(to_unsigned(val, 4));
    end function;

begin

    -- Edge detection process
    process(clk, reset)
        variable T : integer := 0;  -- Declare T variable inside the process
        variable i0, i1, i2, i3 : integer := 0;
        variable F : integer := 0;
    begin
        if reset = '1' then -- clear the output if reset is on
            for i in 0 to 9 loop
                for j in 0 to 9 loop
                    edge_matrix(i, j) <= 0;
                end loop;
            end loop;
        elsif rising_edge(clk) then
            for i in 0 to 9 loop
                for j in 0 to 9 loop
                    edge_matrix(i, j) <= 0;
                end loop;
            end loop;
            -- Calculate the threshold value
            T := compute_threshold(my_matrix);

            -- Iterate over the image matrix to apply edge detection
            for i in 0 to 7 loop  -- count number = no of Rows of the image - no of rows of Gx + 1
                for j in 0 to 7 loop
                    edge_matrix(i, j) <= compute_edge(i, j, T);  
        
                    -- Assertion to check if edge_matrix(i, j) is 1
                    assert edge_matrix(i, j) = 1
                    report "Edge detected at position (" & integer'image(i) & ", " & integer'image(j) & ")" severity note;
                end loop;
            end loop;
            
            -- Find the coordinates of the beginning and the end of the Line detection
            for i in 0 to 7 loop
                for j in 0 to 7 loop
                    if (F = 0) then
                        if (edge_matrix(i, j) = 1) then
                            i0 := i;
                            i1 := j;
                            F  := 1;
                        end if;
                    else  
                        if (edge_matrix(i, j) = 1) then
                            i2 := i;
                            i3 := j;
                        end if;
                    end if;
                end loop;
            end loop;
        end if;

        -- Convert integers to BCD for 7-segment display
        i0_signal <= int_to_bcd(i0);
        i1_signal <= int_to_bcd(i1);
        i2_signal <= int_to_bcd(i2);
        i3_signal <= int_to_bcd(i3);

    end process;

    -- Instantiate 7-segment controllers
    SevenSeg_i0 : entity work.SevenSegmentController
        port map(
            digit => i0_signal,
            segments => segmentsL_i0
        );

    SevenSeg_i1 : entity work.SevenSegmentController
        port map(
            digit => i1_signal,
            segments => segmentsL_i1
        );

    SevenSeg_i2 : entity work.SevenSegmentController
        port map(
            digit => i2_signal,
            segments => segmentsL_i2
        );

    SevenSeg_i3 : entity work.SevenSegmentController
        port map(
            digit => i3_signal,
            segments => segmentsL_i3
        );

end STRUCT;
